**.subckt DAC_10bit_testbench
V8 Vdd GND 1.8
V4 D1 GND pulse 0 1.8 2u .1n .1n 2u 4u
V21 D2 GND pulse 0 1.8 4u .1n .1n 4u 8u
V5 D3 GND pulse 0 1.8 8u .1n .1n 8u 16u
V1 In1 GND 1.8
V2 In2 GND 0
V3 D4 GND pulse 0 1.8 16u .1n .1n 16u 32u
V6 D5 GND pulse 0 1.8 32u .1n .1n 32u 64u
V7 D6 GND pulse 0 1.8 64u .1n .1n 64u 128u
V9 D7 GND pulse 0 1.8 128u .1n .1n 128u 256u
V10 D0 GND pulse 0 1.8 1u .1n .1n 1u 2u
V11 D8 GND pulse 0 1.8 256u .1n .1n 256u 512u
V12 D9 GND pulse 0 1.8 512u .1n .1n 512u 1024u
x1 Vdd out D3 D2 D1 D0 In2 D4 D5 D6 D7 D8 D9 In1 DAC_10bit
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nand3/sky130_fd_sc_hd__nand3_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nand2/sky130_fd_sc_hd__nand2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor3/sky130_fd_sc_hd__nor3_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dfrtp/sky130_fd_sc_hd__dfrtp_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor2/sky130_fd_sc_hd__nor2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dlrbn/sky130_fd_sc_hd__dlrbn_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a31o/sky130_fd_sc_hd__a31o_2.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a222oi/sky130_fd_sc_hd__a222oi_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/or2/sky130_fd_sc_hd__or2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/o221ai/sky130_fd_sc_hd__o221ai_1.spice


**** end user architecture code
**.ends

* expanding   symbol:  DAC_10bit.sym # of pins=14
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_10bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_10bit.sch
.subckt DAC_10bit  Vdd Out D3 D2 D1 D0 In2 D4 D5 D6 D7 D8 D9 In1
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net1 net2 Vdd D9 TG
x1 Vdd net1 D3 D2 D1 D0 vref1 D4 D5 D6 D7 D8 In1 DAC_9bit
x2 Vdd net2 D3 D2 D1 D0 In2 D4 D5 D6 D7 D8 vref1 DAC_9bit
.ends


* expanding   symbol:  TG.sym # of pins=5
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/TG.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/TG.sch
.subckt TG  Out In1 In2 Vdd D
XM1 Dinv D GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 Dinv D Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 Dinv GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net1 Dinv Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 Out net1 In2 In2 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 Out net1 In1 In1 sky130_fd_pr__pfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 In2 Dinv Out Out sky130_fd_pr__pfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 In1 Dinv Out Out sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  DAC_9bit.sym # of pins=13
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_9bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_9bit.sch
.subckt DAC_9bit  Vdd Out D3 D2 D1 D0 In2 D4 D5 D6 D7 D8 In1
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net1 net2 Vdd D8 TG
x1 Vdd net1 D3 D2 D1 D0 vref1 D4 D5 D6 D7 In1 DAC_8bit
x2 Vdd net2 D3 D2 D1 D0 In2 D4 D5 D6 D7 vref1 DAC_8bit
.ends


* expanding   symbol:  DAC_8bit.sym # of pins=12
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_8bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_8bit.sch
.subckt DAC_8bit  Vdd Out D3 D2 D1 D0 In2 D4 D5 D6 D7 In1
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net1 net2 Vdd D7 TG
x1 Vdd net1 D3 D2 D1 D0 vref1 D4 D5 D6 In1 DAC_7bit
x2 Vdd net2 D3 D2 D1 D0 In2 D4 D5 D6 vref1 DAC_7bit
.ends


* expanding   symbol:  DAC_7bit.sym # of pins=11
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_7bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_7bit.sch
.subckt DAC_7bit  Vdd Out D3 D2 D1 D0 In2 D4 D5 D6 In1
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net1 net2 Vdd D6 TG
x1 Vdd net1 D3 D2 D1 D0 vref1 D4 D5 In1 DAC_6bit
x2 Vdd net2 D3 D2 D1 D0 In2 D4 D5 vref1 DAC_6bit
.ends


* expanding   symbol:  DAC_6bit.sym # of pins=10
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_6bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_6bit.sch
.subckt DAC_6bit  Vdd Out D3 D2 D1 D0 In2 D4 D5 In1
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net1 net2 Vdd D5 TG
x1 Vdd net1 D3 D2 D1 D0 vref1 D4 In1 DAC_5bit
x2 Vdd net2 D3 D2 D1 D0 In2 D4 vref1 DAC_5bit
.ends


* expanding   symbol:  DAC_5bit.sym # of pins=9
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_5bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_5bit.sch
.subckt DAC_5bit  Vdd Out D3 D2 D1 D0 In2 D4 In1
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net1 net2 Vdd D4 TG
x1 Vdd net1 D3 D2 D1 D0 vref1 In1 DAC_4bit
x2 Vdd net2 D3 D2 D1 D0 In2 vref1 DAC_4bit
.ends


* expanding   symbol:  DAC_4bit.sym # of pins=8
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_4bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_4bit.sch
.subckt DAC_4bit  Vdd Out D3 D2 D1 D0 In2 In1
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net2 net1 Vdd D3 TG
x1 Vdd net2 In1 D2 D1 D0 vref1 DAC_3bit
x2 Vdd net1 vref1 D2 D1 D0 In2 DAC_3bit
.ends


* expanding   symbol:  DAC_3bit.sym # of pins=7
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_3bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_3bit.sch
.subckt DAC_3bit  Vdd Out In1 D2 D1 D0 In2
x1 Vdd net2 In1 D1 D0 vref1 DAC_2bit
x2 Vdd net1 vref1 D1 D0 In2 DAC_2bit
R8 In1 vref1 250 m=1
R6 vref1 In2 250 m=1
x3 out net2 net1 Vdd D2 TG
.ends


* expanding   symbol:  DAC_2bit.sym # of pins=6
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_2bit.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/DAC_2bit.sch
.subckt DAC_2bit  Vdd Out In1 D1 D0 In2
x1 net1 net3 net4 Vdd D0 TG
x2 net2 net5 In2 Vdd D0 TG
x3 out net1 net2 Vdd D1 TG
R1 In1 net3 500 m=1
R2 net3 net4 500 m=1
R3 net4 net5 500 m=1
R4 net5 In2 500 m=1
.ends

.GLOBAL GND
**** begin user architecture code


.temp 25
vvcc vcc 0 1.8
vvss vss 0 0
.control
tran 1.5m 2048u
plot out
.endc


**** end user architecture code
** flattened .save nodes
.end
