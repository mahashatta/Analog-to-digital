**.subckt stair
V1 A GND pwl 0 0.1 0 0.2 1u 0.2 2u 0.2 2u 0.3 3u 0.3 3u 0.4
**.ends
.GLOBAL GND
**** begin user architecture code


.temp 25
vvcc vcc 0 1.8
vvss vss 0 0
.control
tran 10n 10u
plot A
.endc


**** end user architecture code
** flattened .save nodes
.end
