**.subckt cmpOAI_testbench
V3 B8 GND 0.425
V4 A GND pwl 0 0 12.5u 0 12.5u 0.1 12.5u 0.025 22.5u 0.025 22.5u 0.075 32.5u 0.075 32.5u 0.125 42.5u
+ 0.125 42.5u 0.175 52.5u 0.175 52.5u 0.225 62.5u 0.225 62.5u 0.275 72.5u 0.275 72.5u 0.325 82.5u 0.325
+ 82.5u 0.375 92.5u 0.375 92.5u 0.425 102.5u 0.425 102.5u 0.475 112.5u 0.475 112.5u 0.525 122.5u 0.525
+ 122.5u 0.575 132.5u 0.575 132.5u 0.625 142.5u 0.625 142.5u 0.675 152.5u 0.675 152.5u 0.725 162.5u 0.725
+ 162.5u 0.775 172.5u 0.775 172.5u 0.825 182.5u 0.825 182.5u 0.875 192.5u 0.875 192.5u 0.925 202.5u 0.925
+ 202.5u 0.975
V5 clk GND pulse 0 1.8 5n .1n .1n 1u 2u
V1 B7 GND 0.375
V2 B6 GND 0.325
V6 B5 GND 0.275
V7 B4 GND 0.225
V8 B3 GND 0.175
V9 B2 GND 0.125
V10 B1 GND 0.075
V11 VDD GND 1.8
x1 A B1 Q1 clk VDD GND cmpoaisch
x2 A B2 Q2 clk VDD GND cmpoaisch
x3 A B3 Q3 clk VDD GND cmpoaisch
x4 A B4 Q4 clk VDD GND cmpoaisch
x5 A B5 Q5 clk VDD GND cmpoaisch
x6 A B6 Q6 clk VDD GND cmpoaisch
x7 A B7 Q7 clk VDD GND cmpoaisch
x8 A B8 Q8 clk VDD GND cmpoaisch
x9 A B9 Q9 clk VDD GND cmpoaisch
x10 A B10 Q10 clk VDD GND cmpoaisch
V12 B10 GND 0.525
V13 B9 GND 0.475
V14 B13 GND 0.675
V15 B12 GND 0.625
V16 B11 GND 0.575
V17 B15 GND 0.775
V18 B14 GND 0.725
V19 B17 GND 0.875
V20 B16 GND 0.825
V21 B19 GND 0.975
V22 B18 GND 0.925
x11 A B11 Q11 clk VDD GND cmpoaisch
x12 A B12 Q12 clk VDD GND cmpoaisch
x13 A B13 Q13 clk VDD GND cmpoaisch
x14 A B14 Q14 clk VDD GND cmpoaisch
x15 A B15 Q15 clk VDD GND cmpoaisch
x16 A B16 Q16 clk VDD GND cmpoaisch
x17 A B17 Q17 clk VDD GND cmpoaisch
x18 A B18 Q18 clk VDD GND cmpoaisch
x19 A B19 Q19 clk VDD GND cmpoaisch
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nand3/sky130_fd_sc_hd__nand3_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nand2/sky130_fd_sc_hd__nand2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor3/sky130_fd_sc_hd__nor3_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dfrtp/sky130_fd_sc_hd__dfrtp_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor2/sky130_fd_sc_hd__nor2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dlrbn/sky130_fd_sc_hd__dlrbn_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a31o/sky130_fd_sc_hd__a31o_2.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a222oi/sky130_fd_sc_hd__a222oi_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/or2/sky130_fd_sc_hd__or2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/o221ai/sky130_fd_sc_hd__o221ai_1.spice


**** end user architecture code
**.ends

* expanding   symbol:  cmpoaisch.sym # of pins=6
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/cmpoaisch.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/cmpoaisch.sch
.subckt cmpoaisch  A B Q clk VDD VSS
V7 VNB GND 0
V8 VPWR GND 1.8
V9 VPB GND 1.8
V10 VGND GND 0
x15 clk VGND VNB VPB VPWR clkb sky130_fd_sc_hd__inv_1
x7 A A clkb VPWR net2 VPWR VGND VNB VPB VPWR net1 sky130_fd_sc_hd__a222oi_1
x8 B B clkb VPWR net1 VPWR VGND VNB VPB VPWR net2 sky130_fd_sc_hd__a222oi_1
x10 net1 VGND VNB VPB VPWR net4 sky130_fd_sc_hd__inv_1
x11 net2 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__inv_1
x12 net4 Q VGND VNB VPB VPWR Qd sky130_fd_sc_hd__nand2_1
x13 Qd net3 VGND VNB VPB VPWR Q sky130_fd_sc_hd__nand2_1
.ends

.GLOBAL GND
**** begin user architecture code


.temp 25
vvcc vcc 0 1.8
vvss vss 0 0
.control
tran 0.1u 210u
plot A CLK+2 Q1+4 Q2+6 Q3+8 Q4+10 Q5+12 Q6+14 Q7+16 Q8+18 Q9+20 Q10+22 Q11+24 Q12+26 Q13+28 Q14+30
+ Q15+32 Q16+34 Q17+36 Q18+38 Q19+40
.endc


**** end user architecture code
** flattened .save nodes
.end
