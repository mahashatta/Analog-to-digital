**.subckt cmpoaisch
V7 VNB GND 0
V8 VPWR GND 1.8
V9 VPB GND 1.8
V10 VGND GND 0
x15 clk VGND VNB VPB VPWR clkb sky130_fd_sc_hd__inv_1
x7 A A clkb VPWR net2 VPWR VGND VNB VPB VPWR net1 sky130_fd_sc_hd__a222oi_1
x8 B B clkb VPWR net1 VPWR VGND VNB VPB VPWR net2 sky130_fd_sc_hd__a222oi_1
x10 net1 VGND VNB VPB VPWR net4 sky130_fd_sc_hd__inv_1
x11 net2 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__inv_1
x12 net4 Q VGND VNB VPB VPWR Qd sky130_fd_sc_hd__nand2_1
x13 Qd net3 VGND VNB VPB VPWR Q sky130_fd_sc_hd__nand2_1
**.ends
.GLOBAL GND
** flattened .save nodes
.end
