**.subckt cmpoaisch_2
V7 VNB GND 0
V8 VPWR GND 1.8
V9 VPB GND 1.8
V10 VGND GND 0
x15 clk VGND VNB VPB VPWR clkb sky130_fd_sc_hd__inv_1
x10 net1 VGND VNB VPB VPWR net5 sky130_fd_sc_hd__inv_1
x11 net2 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__inv_1
x1 A A clk GND net2 VGND VNB VPB VPWR net1 sky130_fd_sc_hd__o221a_1
x2 B B clk GND net1 VGND VNB VPB VPWR net2 sky130_fd_sc_hd__o221a_1
x3 net5 Q VGND VNB VPB VPWR net4 sky130_fd_sc_hd__nand2_1
x4 net4 net3 VGND VNB VPB VPWR Q sky130_fd_sc_hd__nand2_1
**.ends
.GLOBAL GND
** flattened .save nodes
.end
