**.subckt cmpoai_all__
x15 clk VGND VNB VPB VPWR clkb sky130_fd_sc_hd__inv_1
x2 net3 VGND VNB VPB VPWR net6 sky130_fd_sc_hd__inv_1
x3 net4 VGND VNB VPB VPWR net5 sky130_fd_sc_hd__inv_1
x6 net4 GND clk GND A VGND VNB VPB VPWR net3 sky130_fd_sc_hd__o221ai_1
x9 net3 GND clk GND B VGND VNB VPB VPWR net4 sky130_fd_sc_hd__o221ai_1
x10 net5 net1 net7 VGND VNB VPB VPWR Q sky130_fd_sc_hd__nor3_1
x11 Q net6 net2 VGND VNB VPB VPWR net7 sky130_fd_sc_hd__nor3_1
x1 A A clkb net2 VGND VNB VPB VPWR net1 sky130_fd_sc_hd__a211oi_1
x4 B B clkb net1 VGND VNB VPB VPWR net2 sky130_fd_sc_hd__a211oi_1
**.ends
.GLOBAL GND
** flattened .save nodes
.end
