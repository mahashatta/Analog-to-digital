**.subckt cmpOAI_all_testbench_
V5 clk GND pulse 0 1.8 2u .1n .1n 2u 4u
V11 VDD GND 1.8
V16 B8 GND 0.7
V17 A1 GND pwl 0 0 12.5u 0 12.5u 0.01 22.5u 0.01 22.5u 0.02 32.5u 0.02 32.5u 0.03 42.5u 0.03 42.5u
+ 0.04 52.5u 0.04 52.5u 0.05 62.5u 0.05 62.5u 0.06 72.5u 0.06 72.5u 0.07 82.5u 0.07 82.5u 0.08 92.5u 0.08
+ 92.5u 0.09 102.5u 0.09 102.5u 0.1 112.5u 0.1
V19 B7 GND 0.6
V20 B6 GND 0.5
V21 B5 GND 0.4
V22 B4 GND 0.3
V23 B3 GND 0.2
V24 B2 GND 0.1
V25 B1 GND 0
V27 B10 GND 0.9
V28 B9 GND 0.8
V30 B12 GND 1.1
V31 B11 GND 1.0
V1 B14 GND 1.3
V2 B13 GND 1.2
V3 B16 GND 1.5
V4 B15 GND 1.4
V6 B18 GND 1.7
V7 B17 GND 1.6
V8 A2 GND pwl 0 0.1 12.5u 0.1 12.5u 0.11 22.5u 0.11 22.5u 0.12 32.5u 0.12 32.5u 0.13 42.5u 0.13
+ 42.5u 0.14 52.5u 0.14 52.5u 0.15 62.5u 0.15 62.5u 0.16 72.5u 0.16 72.5u 0.17 82.5u 0.17 82.5u 0.18 92.5u
+ 0.18 92.5u 0.19 102.5u 0.19 102.5u 0.2 112.5u 0.2
V9 A3 GND pwl 0 0.2 12.5u 0.2 12.5u 0.21 22.5u 0.21 22.5u 0.22 32.5u 0.22 32.5u 0.23 42.5u 0.23
+ 42.5u 0.24 52.5u 0.24 52.5u 0.25 62.5u 0.25 62.5u 0.26 72.5u 0.26 72.5u 0.27 82.5u 0.27 82.5u 0.28 92.5u
+ 0.28 92.5u 0.29 102.5u 0.29 102.5u 0.3 112.5u 0.3
V10 A4 GND pwl 0 0.3 12.5u 0.3 12.5u 0.31 22.5u 0.31 22.5u 0.32 32.5u 0.32 32.5u 0.33 42.5u 0.33
+ 42.5u 0.34 52.5u 0.34 52.5u 0.35 62.5u 0.35 62.5u 0.36 72.5u 0.36 72.5u 0.37 82.5u 0.37 82.5u 0.38 92.5u
+ 0.38 92.5u 0.39 102.5u 0.39 102.5u 0.4 112.5u 0.4
V12 A5 GND pwl 0 0.4 12.5u 0.4 12.5u 0.41 22.5u 0.41 22.5u 0.42 32.5u 0.42 32.5u 0.43 42.5u 0.43
+ 42.5u 0.44 52.5u 0.44 52.5u 0.45 62.5u 0.45 62.5u 0.46 72.5u 0.46 72.5u 0.47 82.5u 0.47 82.5u 0.48 92.5u
+ 0.48 92.5u 0.49 102.5u 0.49 102.5u 0.5 112.5u 0.5
V13 A6 GND pwl 0 0.5 12.5u 0.5 12.5u 0.51 22.5u 0.51 22.5u 0.52 32.5u 0.52 32.5u 0.53 42.5u 0.53
+ 42.5u 0.54 52.5u 0.54 52.5u 0.55 62.5u 0.55 62.5u 0.56 72.5u 0.56 72.5u 0.57 82.5u 0.57 82.5u 0.58 92.5u
+ 0.58 92.5u 0.59 102.5u 0.59 102.5u 0.6 112.5u 0.6
V14 A7 GND pwl 0 0.6 12.5u 0.6 12.5u 0.61 22.5u 0.61 22.5u 0.62 32.5u 0.62 32.5u 0.63 42.5u 0.63
+ 42.5u 0.64 52.5u 0.64 52.5u 0.65 62.5u 0.65 62.5u 0.66 72.5u 0.66 72.5u 0.67 82.5u 0.67 82.5u 0.68 92.5u
+ 0.68 92.5u 0.69 102.5u 0.69 102.5u 0.7 112.5u 0.7
V15 A8 GND pwl 0 0.7 12.5u 0.7 12.5u 0.71 22.5u 0.71 22.5u 0.72 32.5u 0.72 32.5u 0.73 42.5u 0.73
+ 42.5u 0.74 52.5u 0.74 52.5u 0.75 62.5u 0.75 62.5u 0.76 72.5u 0.76 72.5u 0.77 82.5u 0.77 82.5u 0.78 92.5u
+ 0.78 92.5u 0.79 102.5u 0.79 102.5u 0.8 112.5u 0.8
V18 A9 GND pwl 0 .8 12.5u 0.8 12.5u 0.81 22.5u 0.81 22.5u 0.82 32.5u 0.82 32.5u 0.83 42.5u 0.83
+ 42.5u 0.84 52.5u 0.84 52.5u 0.85 62.5u 0.85 62.5u 0.86 72.5u 0.86 72.5u 0.87 82.5u 0.87 82.5u 0.88 92.5u
+ 0.88 92.5u 0.89 102.5u 0.89 102.5u 0.9 112.5u 0.9
V26 A10 GND pwl 0 0.9 12.5u 0.9 12.5u 0.91 22.5u 0.91 22.5u 0.92 32.5u 0.92 32.5u 0.93 42.5u 0.93
+ 42.5u 0.94 52.5u 0.94 52.5u 0.95 62.5u 0.95 62.5u 0.96 72.5u 0.96 72.5u 0.97 82.5u 0.97 82.5u 0.98 92.5u
+ 0.98 92.5u 0.99 102.5u 0.99 102.5u 1.0 112.5u 1.0
V29 A11 GND pwl 0 1.0 12.5u 1.0 12.5u 1.01 22.5u 1.01 22.5u 1.02 32.5u 1.02 32.5u 1.03 42.5u 1.03
+ 42.5u 1.04 52.5u 1.04 52.5u 1.05 62.5u 1.05 62.5u 1.06 72.5u 1.06 72.5u 1.07 82.5u 1.07 82.5u 1.08 92.5u
+ 1.08 92.5u 1.09 102.5u 1.09 102.5u 1.1 112.5u 1.1
V32 A12 GND pwl 0 1.1 12.5u 1.1 12.5u 1.11 22.5u 1.11 22.5u 1.12 32.5u 1.12 32.5u 1.13 42.5u 1.13
+ 42.5u 1.14 52.5u 1.14 52.5u 1.15 62.5u 1.15 62.5u 1.16 72.5u 1.16 72.5u 1.17 82.5u 1.17 82.5u 1.18 92.5u
+ 1.18 92.5u 1.19 102.5u 1.19 102.5u 1.2 112.5u 1.2
V33 A13 GND pwl 0 1.2 12.5u 1.2 12.5u 1.21 22.5u 1.21 22.5u 1.22 32.5u 1.22 32.5u 1.23 42.5u 1.23
+ 42.5u 1.24 52.5u 1.24 52.5u 1.25 62.5u 1.25 62.5u 1.26 72.5u 1.26 72.5u 1.27 82.5u 1.27 82.5u 1.28 92.5u
+ 1.28 92.5u 1.29 102.5u 1.29 102.5u 1.3 112.5u 1.3
V34 A14 GND pwl 0 1.3 12.5u 1.3 12.5u 1.31 22.5u 1.31 22.5u 1.32 32.5u 1.32 32.5u 1.33 42.5u 1.33
+ 42.5u 1.34 52.5u 1.34 52.5u 1.35 62.5u 1.35 62.5u 1.36 72.5u 1.36 72.5u 1.37 82.5u 1.37 82.5u 1.38 92.5u
+ 1.38 92.5u 1.39 102.5u 1.39 102.5u 1.4 112.5u 1.4
V35 A15 GND pwl 0 1.4 12.5u 1.4 12.5u 1.41 22.5u 1.41 22.5u 1.42 32.5u 1.42 32.5u 1.43 42.5u 1.43
+ 42.5u 1.44 52.5u 1.44 52.5u 1.45 62.5u 1.45 62.5u 1.46 72.5u 1.46 72.5u 1.47 82.5u 1.47 82.5u 1.48 92.5u
+ 1.48 92.5u 1.49 102.5u 1.49 102.5u 1.5 112.5u 1.5
V36 A16 GND pwl 0 1.5 12.5u 1.5 12.5u 1.51 22.5u 1.51 22.5u 1.52 32.5u 1.52 32.5u 1.53 42.5u 1.53
+ 42.5u 1.54 52.5u 1.54 52.5u 1.55 62.5u 1.55 62.5u 1.56 72.5u 1.56 72.5u 1.57 82.5u 1.57 82.5u 1.58 92.5u
+ 1.58 92.5u 1.59 102.5u 1.59 102.5u 1.6 112.5u 1.6
V37 A17 GND pwl 0 1.6 12.5u 1.6 12.5u 1.61 22.5u 1.61 22.5u 1.62 32.5u 1.62 32.5u 1.63 42.5u 1.63
+ 42.5u 1.64 52.5u 1.64 52.5u 1.65 62.5u 1.65 62.5u 1.66 72.5u 1.66 72.5u 1.67 82.5u 1.67 82.5u 1.68 92.5u
+ 1.68 92.5u 1.69 102.5u 1.69 102.5u 1.7 112.5u 1.7
V38 A18 GND pwl 0 1.7 12.5u 1.7 12.5u 1.71 22.5u 1.71 22.5u 1.72 32.5u 1.72 32.5u 1.73 42.5u 1.73
+ 42.5u 1.74 52.5u 1.74 52.5u 1.75 62.5u 1.75 62.5u 1.76 72.5u 1.76 72.5u 1.77 82.5u 1.77 82.5u 1.78 92.5u
+ 1.78 92.5u 1.79 102.5u 1.79 102.5u 1.8 112.5u 1.8
x1 A1 B1 Q1 clk VDD GND VDD GND cmpoai_all__
x2 A2 B2 Q2 clk VDD GND VDD GND cmpoai_all__
x3 A3 B3 Q3 clk VDD GND VDD GND cmpoai_all__
x4 A4 B4 Q4 clk VDD GND VDD GND cmpoai_all__
x5 A5 B5 Q5 clk VDD GND VDD GND cmpoai_all__
x6 A6 B6 Q6 clk VDD GND VDD GND cmpoai_all__
x7 A7 B7 Q7 clk VDD GND VDD GND cmpoai_all__
x8 A8 B8 Q8 clk VDD GND VDD GND cmpoai_all__
x9 A9 B9 Q9 clk VDD GND VDD GND cmpoai_all__
x10 A10 B10 Q10 clk VDD GND VDD GND cmpoai_all__
x11 A11 B11 Q11 clk VDD GND VDD GND cmpoai_all__
x12 A12 B12 Q12 clk VDD GND VDD GND cmpoai_all__
x13 A13 B13 Q13 clk VDD GND VDD GND cmpoai_all__
x14 A14 B14 Q14 clk VDD GND VDD GND cmpoai_all__
x15 A15 B15 Q15 clk VDD GND VDD GND cmpoai_all__
x16 A16 B16 Q16 clk VDD GND VDD GND cmpoai_all__
x17 A17 B17 Q17 clk VDD GND VDD GND cmpoai_all__
x18 A18 B18 Q18 clk VDD GND VDD GND cmpoai_all__
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nand3/sky130_fd_sc_hd__nand3_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nand2/sky130_fd_sc_hd__nand2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor3/sky130_fd_sc_hd__nor3_4.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor3/sky130_fd_sc_hd__nor3_2.spice

.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor3/sky130_fd_sc_hd__nor3_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dfrtp/sky130_fd_sc_hd__dfrtp_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/nor2/sky130_fd_sc_hd__nor2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dlrbn/sky130_fd_sc_hd__dlrbn_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a31o/sky130_fd_sc_hd__a31o_2.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_2.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a222oi/sky130_fd_sc_hd__a222oi_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a221oi/sky130_fd_sc_hd__a221oi_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/a221oi/sky130_fd_sc_hd__a221oi_4.spice

.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/or2/sky130_fd_sc_hd__or2_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/o221ai/sky130_fd_sc_hd__o221ai_1.spice
.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/o221ai/sky130_fd_sc_hd__o221ai_4.spice



**** end user architecture code
**.ends

* expanding   symbol:  cmpoai_all__.sym # of pins=8
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/cmpoai_all__.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/cmpoai_all__.sch
.subckt cmpoai_all__  A B Q clk VPB VNB VPWR VGND
x15 clk VGND VNB VPB VPWR clkb sky130_fd_sc_hd__inv_1
x7 VPWR net2 clkb VPWR A VGND VNB VPB VPWR net1 sky130_fd_sc_hd__a221oi_1
x8 net1 VPWR clkb VPWR B VGND VNB VPB VPWR net2 sky130_fd_sc_hd__a221oi_1
x2 net3 VGND VNB VPB VPWR net6 sky130_fd_sc_hd__inv_1
x3 net4 VGND VNB VPB VPWR net5 sky130_fd_sc_hd__inv_1
x6 net4 GND clk GND A VGND VNB VPB VPWR net3 sky130_fd_sc_hd__o221ai_1
x9 net3 GND clk GND B VGND VNB VPB VPWR net4 sky130_fd_sc_hd__o221ai_1
x10 net5 net1 net7 VGND VNB VPB VPWR Q sky130_fd_sc_hd__nor3_1
x11 Q net6 net2 VGND VNB VPB VPWR net7 sky130_fd_sc_hd__nor3_1
.ends

.GLOBAL GND
**** begin user architecture code


.temp 25
vvcc vcc 0 1.8
vvss vss 0 0
.control
tran 0.5u 130u
plot Q1 Q2+2 Q3+4 Q4+6 Q5+8 Q6+10 Q7+12 Q8+14 Q9+16 Q10+18 Q11+20 Q12+22 Q13+24 Q14+28 Q15+30 Q16+32
+ Q17+34 Q18+36
meas tran x find t(Q1) when v(Q1)=1.8
meas tran x find t(Q2) when v(Q2)=1.8
meas tran x find t(Q3) when v(Q3)=1.8
meas tran x find t(Q4) when v(Q4)=1.8
meas tran x find t(Q5) when v(Q5)=1.8
meas tran x find t(Q6) when v(Q6)=1.8
meas tran x find t(Q7) when v(Q7)=1.8
meas tran x find t(Q8) when v(Q8)=1.8
meas tran x find t(Q9) when v(Q9)=1.8
meas tran x find t(Q10) when v(Q10)=1.8
meas tran x find t(Q11) when v(Q11)=1.8
meas tran x find t(Q12) when v(Q12)=1.8
meas tran x find t(Q13) when v(Q13)=1.8
meas tran x find t(Q14) when v(Q14)=1.8
meas tran x find t(Q15) when v(Q15)=1.8
meas tran x find t(Q16) when v(Q16)=1.8
meas tran x find t(Q17) when v(Q17)=1.8
meas tran x find t(Q18) when v(Q18)=1.8

.endc


**** end user architecture code
** flattened .save nodes
.end
