**.subckt test_comparator CAL PLUS MINUS EN VSS VCC SAOUT
*.ipin CAL
*.ipin PLUS
*.ipin MINUS
*.ipin EN
*.ipin VSS
*.ipin VCC
*.opin SAOUT
E5 TEMPERAT VSS VOL=' temper ' 
C38 VSS 0 2p m=1
C3 SAOUTF 0 4f m=1
C5 GN 0 4f m=1
C30 SN 0 2f m=1
C31 OUTDIFF 0 4f m=1
v2 net1 VSSI 0
v3 net4 VSSI 0
v4 net3 VSSI 0
v6 net2 VSSI 0
C1 SAOUT 0 4f m=1
v1 net5 VSSI 0
v5 net6 VSSI 0
C7 GP 0 4f m=1
x4 CALBB CALB VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x5 CALB CAL VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
XM4 SP VSS VCC VCC sky130_fd_pr__pfet_01v8 L=1 W=0.55 nf=1 ad='W * 0.29' as='W * 0.29' pd='W + 2 * 0.29'
+ ps='W + 2 * 0.29' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM5 OUTDIFF GN VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM6 GN GN VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM8 SAOUTF OUTDIFF VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM9 SAOUT SAOUTF VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM11 SAOUT EN VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='W + 2 * 0.29'
+ ps='W + 2 * 0.29' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM12 SAOUT ZERO2 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=0.42 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM13 SAOUTF ZERO1 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=0.42 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM14 OUTDIFF ZERO0 VCC VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=0.42 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM1 VSSI EN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='W + 2 * 0.29'
+ ps='W + 2 * 0.29' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=2 m=2 
XM2 OUTDIFF ZERO0 net2 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=0.42 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM3 SAOUTF ZERO1 net3 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=0.42 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM7 SAOUT ZERO2 net6 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=0.42 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM15 SAOUT SAOUTF net5 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM10 SAOUTF OUTDIFF net4 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM17 SN VCC net1 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=0.42 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM18 OUTDIFF GP VSSI VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM19 GP GP VSSI VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM20 OUTDIFF PLUS SP VCC sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM21 GP MINUS SP VCC sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM23 OUTDIFF PLUS SN VSS sky130_fd_pr__nfet_01v8_lvt L=0.25 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
XM16 GN MINUS SN VSS sky130_fd_pr__nfet_01v8_lvt L=0.25 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1 
x1 OUTDIFF ZERO0 CALB CALBB VCC VSS passgate_nlvt W_N=0.42 L_N=0.15 W_P=0.42 L_P=0.15 m=1
x2 SAOUTF ZERO1 CALB CALBB VCC VSS passgate_nlvt W_N=0.42 L_N=0.15 W_P=0.42 L_P=0.15 m=1
x3 SAOUT ZERO2 CALB CALBB VCC VSS passgate_nlvt W_N=0.42 L_N=0.15 W_P=0.42 L_P=0.15 m=1
C2 ZERO0 VCC 15f m=1
C4 ZERO1 VCC 15f m=1
C6 ZERO2 VCC 15f m=1
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice

**** end user architecture code
**.ends

* expanding   symbol:  sky130_tests/not.sym # of pins=2
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/sky130_tests/not.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/sky130_tests/not.sch
.subckt not  y a  VCCPIN  VSSPIN      W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sky130_tests/passgate_nlvt.sym # of pins=4
* sym_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/sky130_tests/passgate_nlvt.sym
* sch_path: /home/mahashatta/.xschem/xschem_library/xschem_sky130/sky130_tests/passgate_nlvt.sch
.subckt passgate_nlvt  Z A GP GN  VCCBPIN  VSSBPIN   W_N=1 L_N=0.35 W_P=1 L_P=0.35
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8_lvt L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8_lvt L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

**** begin user architecture code

* .option SCALE=1e-6
.option method=gear seed=12

* this experimental option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1

* .param VCC=1.8
.param VCCGAUSS=agauss(1.8, 0.05, 1)
.param VCC=VCCGAUSS
.param VDL='VCC/2+0.2'
.param ABSVAR=0.02
.temp 25

** to generate following file:
** copy .../xschem_sky130/sky130_tests/stimuli.test_comparator to simulation directory
** then do 'Simulation->Utile Stimuli Editor (GUI)' and press 'Translate'
.include "stimuli_test_comparator.cir"

** variation marameters:
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre='agauss(0, ABSVAR, 3)/sky130_fd_pr__nfet_01v8_lvt__vth0_slope'
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre='agauss(0, ABSVAR, 3)/sky130_fd_pr__pfet_01v8_lvt__vth0_slope'

* .tran 0.1n 900n uic

.control
  let run=1
  dowhile run <= 20
    if run > 1
      reset
      set appendwrite
    end
    save all
    * save saout cal i(vvcc) en plus minus
    tran 0.1n 300n uic
    write test_comparator.raw
    let run = run + 1
  end
.endc


**** end user architecture code
** flattened .save nodes
.save I(v2)
.save I(v3)
.save I(v4)
.save I(v6)
.save I(v1)
.save I(v5)
.end
